`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/10/23 14:11:51
// Design Name: 
// Module Name: prng_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module prng_top(
    clk,
    rstn,
    data_out,
    get_random
    );

/////////////////////////////////////////////////////////////////////////////////
//  I/O
/////////////////////////////////////////////////////////////////////////////////
input               clk;
input               rstn;
input               get_random;

output      [7:0]   data_out;

/////////////////////////////////////////////////////////////////////////////////
// def 
/////////////////////////////////////////////////////////////////////////////////
parameter   seed = 32'h02468acd;
wire        [31:0]  lfsr;
wire                data_done;
wire        [1:0]   cnt;

/////////////////////////////////////////////////////////////////////////////////
// fsm 
/////////////////////////////////////////////////////////////////////////////////
assign      data_done = cnt == 2'b11;   
wire        [1:0]   state;

parameter   IDLE = 2'b00;
parameter   SHIFT = 2'b01;
parameter   DATAOUT = 2'b10;
wire        state_shift = state == SHIFT;
wire        state_dataout = state == DATAOUT;

fsm _fsm(
    .clk            (clk            ),
    .rstn           (rstn           ),
    .data_done      (data_done      ),
    .get_random     (get_random     ),
    .state          (state          )
);


/////////////////////////////////////////////////////////////////////////////////
// lfsr 
/////////////////////////////////////////////////////////////////////////////////
prng_lfsr _prng_lfsr(
    .clk            (clk            ),
    .rstn           (rstn           ),
    .seed_load      (1'b0           ),
    .seed           (seed           ),
    .shift_en       (state_shift    ),
    .lfsr           (lfsr           )
);

/////////////////////////////////////////////////////////////////////////////////
// counter 
/////////////////////////////////////////////////////////////////////////////////
prng_counter _prng_counter(
    .clk            (clk            ),   
    .rstn           (rstn           ),
    .cnt_en         (state_dataout  ),
    .cnt            (cnt            )
);

/////////////////////////////////////////////////////////////////////////////////
// output 
/////////////////////////////////////////////////////////////////////////////////
assign data_out = state_dataout ? lfsr >> {cnt,3'b0} : 8'b0;


endmodule
